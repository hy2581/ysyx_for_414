module EXU (
    input clk,
    input rst,
    input [31:0] op,      
    input op_en,          // 只会置于1一周期
    input [31:0] pc,      // 当前指令的PC
    
    output reg ex_end,    // 在处理结束时使得ex_end=!ex_end
    output reg [31:0] next_pc, // 下一条指令的PC
    output reg branch_taken,   // 分支是否taken
    output reg ebreak_flag,     // ebreak 指令执行标志
    output reg [31:0] exit_code, // 添加退出码输出
    
    // 内存接口
    output reg mem_read,       // 内存读使能
    output reg mem_write,      // 内存写使能
    output reg [31:0] mem_addr, // 内存地址
    output reg [31:0] mem_wdata, // 写入内存的数据
    output reg [3:0] mem_mask,   // 字节使能
    input [31:0] mem_rdata,      // 从内存读取的数据
    
    // 添加寄存器接口用于DiffTest
    output [31:0] regs [0:31]
);
    
    // 定义寄存器和信号
    reg [31:0] wdata;
    reg [4:0] waddr;  
    reg wen;//write_en
    reg [4:0] raddr1;
    reg [4:0] raddr2;
    wire [31:0] rdata1;
    wire [31:0] rdata2;
    
    // 操作码和功能码提取
    wire [6:0] opcode = op[6:0];
    wire [2:0] funct3 = op[14:12];
    wire [6:0] funct7 = op[31:25];
    wire [4:0] rd = op[11:7];     // 目标寄存器
    wire [4:0] rs1 = op[19:15];   // 源寄存器1
    wire [4:0] rs2 = op[24:20];   // 源寄存器2
    
    // 各类型立即数解码
    wire [11:0] imm_i = op[31:20];                      // I型立即数
    wire [11:0] imm_s = {op[31:25], op[11:7]};          // S型立即数
    wire [12:0] imm_b = {op[31], op[7], op[30:25], op[11:8], 1'b0}; // B型立即数
    wire [31:0] imm_u = {op[31:12], 12'b0};             // U型立即数
    wire [20:0] imm_j = {op[31], op[19:12], op[20], op[30:21], 1'b0}; // J型立即数
    
    // 扩展后的立即数
    wire [31:0] imm_i_sext = {{20{imm_i[11]}}, imm_i};
    wire [31:0] imm_s_sext = {{20{imm_s[11]}}, imm_s};
    wire [31:0] imm_b_sext = {{19{imm_b[12]}}, imm_b};
    wire [31:0] imm_j_sext = {{11{imm_j[20]}}, imm_j};
    
    // 指令状态
    reg [2:0] state;
    parameter IDLE = 3'b000;
    parameter DECODE = 3'b001;
    parameter EXECUTE = 3'b010;
    parameter MEMORY = 3'b011;
    parameter WRITEBACK = 3'b100;

    // 组合分支条件（避免在时序块里先非阻塞赋值再使用造成时序问题）
    wire branch_cond = (funct3 == 3'b000) ? (rdata1 == rdata2) :
                       (funct3 == 3'b001) ? (rdata1 != rdata2) :
                       (funct3 == 3'b100) ? ($signed(rdata1) < $signed(rdata2)) :
                       (funct3 == 3'b101) ? ($signed(rdata1) >= $signed(rdata2)) :
                       (funct3 == 3'b110) ? (rdata1 < rdata2) :
                       (funct3 == 3'b111) ? (rdata1 >= rdata2) :
                       1'b0;
    
    // 修改寄存器状态检查方法
    // 由于无法直接访问i0.regs，我们使用32个单独的wire来获取寄存器值
    wire [31:0] reg_values [0:31];
    
    // 修改后的寄存器文件实例化，添加寄存器值输出
    RegisterFile #(.ADDR_WIDTH(5), .DATA_WIDTH(32)) i0 (
        .clk(clk),
        .rst(rst),
        .wdata(wdata),
        .waddr(waddr),
        .wen(wen),
        .raddr1(raddr1),
        .rdata1(rdata1),
        .raddr2(raddr2),
        .rdata2(rdata2),
        .reg_values(reg_values)  // 添加这一行用于获取所有寄存器值
    );
    
    // 内存访问临时存储
    reg [31:0] mem_result;
    
    // 指令执行状态机
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= IDLE;
            ex_end <= 0;
            wen <= 0;
            branch_taken <= 0;
            next_pc <= 0;
            mem_read <= 0;
            mem_write <= 0;
            ebreak_flag <= 0;
        end else begin
            case (state)
                IDLE: begin
                    if (op_en) begin
                        state <= DECODE;
                        wen <= 0;
                        branch_taken <= 0;
                        
                        mem_read <= 0;
                        mem_write <= 0;
                        ebreak_flag <= 0;  // 清除 ebreak 标志
                    end
                end
                
                DECODE: begin
                    // 其实没必要，这里强行多打了一拍
                    raddr1 <= rs1[4:0]; 
                    raddr2 <= rs2[4:0];
                    state <= EXECUTE;
                end
                
                EXECUTE: begin
                    case (opcode)
                        // R型指令 - 寄存器-寄存器运算
                        7'b0110011: begin
                            waddr <= rd[4:0];
                            wen <= 1;
                            next_pc <= pc + 4; // 默认PC+4
                            
                            case ({funct7, funct3})
                                // ADD
                                10'b0000000_000: wdata <= rdata1 + rdata2;
                                // SUB
                                10'b0100000_000: wdata <= rdata1 - rdata2;
                                // SLL
                                10'b0000000_001: wdata <= rdata1 << rdata2[4:0];
                                // SLT
                                10'b0000000_010: wdata <= ($signed(rdata1) < $signed(rdata2)) ? 32'b1 : 32'b0;
                                // SLTU
                                10'b0000000_011: wdata <= (rdata1 < rdata2) ? 32'b1 : 32'b0;
                                // XOR
                                10'b0000000_100: wdata <= rdata1 ^ rdata2;
                                // SRL
                                10'b0000000_101: wdata <= rdata1 >> rdata2[4:0];
                                // SRA
                                10'b0100000_101: wdata <= $signed(rdata1) >>> rdata2[4:0];
                                // OR
                                10'b0000000_110: wdata <= rdata1 | rdata2;
                                // AND
                                10'b0000000_111: wdata <= rdata1 & rdata2;
                                default: wen <= 0;
                            endcase
                            state <= WRITEBACK;
                        end
                        
                        // I型指令 - 立即数运算
                        7'b0010011: begin
                            waddr <= rd[4:0];
                            wen <= 1;
                            next_pc <= pc + 4; // 默认PC+4
                            case (funct3)
                                // ADDI
                                3'b000: wdata <= rdata1 + imm_i_sext;
                                // SLTI
                                3'b010: wdata <= ($signed(rdata1) < $signed(imm_i_sext)) ? 32'b1 : 32'b0;
                                // SLTIU
                                3'b011: wdata <= (rdata1 < imm_i_sext) ? 32'b1 : 32'b0;
                                // XORI
                                3'b100: wdata <= rdata1 ^ imm_i_sext;
                                // ORI
                                3'b110: wdata <= rdata1 | imm_i_sext;
                                // ANDI
                                3'b111: wdata <= rdata1 & imm_i_sext;
                                // SLLI
                                3'b001: wdata <= rdata1 << imm_i[4:0];
                                // SRLI/SRAI
                                3'b101: begin
                                    if (imm_i[11:5] == 7'b0000000)
                                        wdata <= rdata1 >> imm_i[4:0]; // SRLI
                                    else if (imm_i[11:5] == 7'b0100000)
                                        wdata <= $signed(rdata1) >>> imm_i[4:0]; // SRAI
                                    else
                                        wen <= 0;
                                end
                                default: wen <= 0;
                            endcase
                            state <= WRITEBACK;
                        end
                        
                        // 加载指令
                        7'b0000011: begin
                            mem_addr <= rdata1 + imm_i_sext;
                            mem_read <= 1;
                            waddr <= rd[4:0];
                            wen <= 1;
                            next_pc <= pc + 4; // 默认PC+4
                            case (funct3)
                                // LB, LH, LW, LBU, LHU
                                3'b000: mem_mask <= 4'b0001; // LB
                                3'b001: mem_mask <= 4'b0011; // LH
                                3'b010: mem_mask <= 4'b1111; // LW
                                3'b100: mem_mask <= 4'b0001; // LBU
                                3'b101: mem_mask <= 4'b0011; // LHU
                                default: begin
                                    mem_read <= 0;
                                    wen <= 0;
                                end
                            endcase
                            state <= MEMORY;
                        end
                        
                        // 存储指令
                        7'b0100011: begin
                            mem_addr <= rdata1 + imm_s_sext;
                            mem_wdata <= rdata2;
                            mem_write <= 1;
                            next_pc <= pc + 4; // 默认PC+4
                            case (funct3)
                                // SB: 写入从 mem_addr 起始的1字节
                                3'b000: mem_mask <= 4'b0001;
                                // SH: 写入从 mem_addr 起始的2字节（允许非对齐）
                                3'b001: mem_mask <= 4'b0011;
                                // SW: 写入从 mem_addr 起始的4字节（允许非对齐）
                                3'b010: mem_mask <= 4'b1111;
                                default: mem_write <= 0;
                            endcase
                            state <= MEMORY;
                        end
                        
                        // 分支指令
                        7'b1100011: begin
                            // 使用组合信号 branch_cond 计算分支结果，避免 non-blocking 更新顺序问题
                            branch_taken <= branch_cond;
                            // imm_b_sext 已按 B 型立即数符号扩展
                            next_pc <= branch_cond ? (pc + imm_b_sext) : (pc + 4);

                            state <= WRITEBACK;
                        end
                        
                        // JAL
                        7'b1101111: begin
                            waddr <= rd[4:0];
                            wdata <= pc + 4;
                            wen <= 1;
                            next_pc <= pc + imm_j_sext;
                            branch_taken <= 1;
                            state <= WRITEBACK;
                        end
                        
                        // JALR
                        7'b1100111: begin
                            if (funct3 == 3'b000) begin
                                waddr <= rd[4:0];
                                wdata <= pc + 4;
                                wen <= 1;
                                next_pc <= (rdata1 + imm_i_sext) & 32'hFFFFFFFE;
                                branch_taken <= 1;
                            end
                            state <= WRITEBACK;
                        end
                        
                        // LUI
                        7'b0110111: begin
                            waddr <= rd[4:0];
                            wdata <= imm_u;
                            wen <= 1;
                            state <= WRITEBACK;
                            next_pc <= pc + 4; // 默认PC+4
                        end
                        
                        // AUIPC
                        7'b0010111: begin
                            waddr <= rd[4:0];
                            wdata <= pc + imm_u;
                            wen <= 1;
                            state <= WRITEBACK;
                            next_pc <= pc + 4; // 默认PC+4
                        end
                        
                        // SYSTEM 指令 (包含 ebreak)
                        7'b1110011: begin
                            if (funct3 == 3'b000 && imm_i == 12'h001) begin
                                ebreak_flag <= 1;
                                exit_code <= reg_values[10];
                            end
                            next_pc <= pc + 4; // 默认PC+4
                            state <= WRITEBACK;
                        end
                        
                        default: begin
                            wen <= 0;
                            state <= WRITEBACK;
                        end
                    endcase
                    
                end
                
                MEMORY: begin
                    mem_read <= 0;
                    mem_write <= 0;
                    
                    if (opcode == 7'b0000011) begin // 加载指令
                        case (funct3)
                            // LB: 从 mem_addr 起始位置取1字节并符号扩展
                            3'b000: begin
                                wdata <= {{24{mem_rdata[7]}}, mem_rdata[7:0]};
                            end
                            // LH: 从 mem_addr 起始位置取2字节并符号扩展（允许非对齐）
                            3'b001: begin
                                wdata <= {{16{mem_rdata[15]}}, mem_rdata[15:0]};
                            end
                            // LW: 从 mem_addr 起始位置取4字节（允许非对齐）
                            3'b010: begin
                                wdata <= mem_rdata;
                            end
                            // LBU: 从 mem_addr 起始位置取1字节零扩展
                            3'b100: begin
                                wdata <= {24'b0, mem_rdata[7:0]};
                            end
                            // LHU: 从 mem_addr 起始位置取2字节零扩展（允许非对齐）
                            3'b101: begin
                                wdata <= {16'b0, mem_rdata[15:0]};
                            end
                            default: wen <= 0;
                        endcase
                    end
                    
                    state <= WRITEBACK;
                end
                
                WRITEBACK: begin
                    // $display("next_pc=0x%x",next_pc);
                    state <= IDLE;
                    ex_end <= ~ex_end;  // 指令执行完成，切换ex_end信号
                    wen <= 0;
                end
                
                default: state <= IDLE;
            endcase
        end
    end
    
    // 替换有问题的generate块
    genvar i;
    generate
        for (i = 0; i < 32; i = i + 1) begin : REG_OUTPUT
            assign regs[i] = (i == 0) ? 32'b0 : reg_values[i]; // x0永远为0
        end
    endgenerate
    
endmodule